module MyMux
( input test
);
  
endmodule